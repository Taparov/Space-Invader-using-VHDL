--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Num_Txt_Sprite is

-- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
--
-- Declare constants
--
-- constant <constant_name>		: time := <time_unit> ns;
-- constant <constant_name>		: integer := <value;
--
-- Declare functions and procedure
--
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--
	type num_array is array(0 to 9) of std_logic_vector(15 downto 0);
	type sprite_array is array(0 to 9) of num_array;
	type alphabet_array is array(0 to 14) of std_logic_vector(23 downto 0);
	type txt_arr is array (natural range <>) of alphabet_array;
	
	-- Declare a constant sprite array for numbers 0-9
  constant num_sprites : sprite_array := (
    -- Sprite for '0'
    ("0000111111110000",
	  "0000111111110000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000000000000000",
	  "0000000000000000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000111111110000",
	  "0000111111110000"),
    
    -- Sprite for '1'
    ("0000000000000000",
     "0000000000000000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000000000000000",
	  "0000000000000000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000000000000000",
	  "0000000000000000"),

    -- Sprite for '2'
    ("0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000111111110000",
	  "0000111111110000",
	  "0111000000000000",
	  "0111000000000000",
	  "0000111111110000",
	  "0000111111110000"),

    -- Sprite for '3'
    ("0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000111111110000",
	  "0000111111110000"),

    -- Sprite for '4'
    ("0000000000000000",
     "0000000000000000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000000000000000",
     "0000000000000000"),

    -- Sprite for '5'
    ("0000111111110000",
	  "0000111111110000",
	  "0111000000000000",
	  "0111000000000000",
	  "0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000111111110000",
	  "0000111111110000"),

    -- Sprite for '6'
    ("0000111111110000",
	  "0000111111110000",
	  "0111000000000000",
	  "0111000000000000",
	  "0000111111110000",
	  "0000111111110000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000111111110000",
	  "0000111111110000"),

    -- Sprite for '7'
    ("0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000000000000000",
	  "0000000000000000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000000000000000",
	  "0000000000000000"),

    -- Sprite for '8'
    ("0000111111110000",
	  "0000111111110000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000111111110000",
	  "0000111111110000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000111111110000",
	  "0000111111110000"),

    -- Sprite for '9'
    ("0000111111110000",
	  "0000111111110000",
	  "0111000000001110",
	  "0111000000001110",
	  "0000111111110000",
	  "0000111111110000",
	  "0000000000001110",
	  "0000000000001110",
	  "0000111111110000",
	  "0000111111110000")
  );
  
  constant game_over_spt : txt_arr (0 to 3) := (
	("001111110000000000000000",
	 "001111111110000000000000",
	 "001110000001110000000000",
	 "001110000000001110000000",
	 "001110000000000111100000",
	 "001110000000000000111000",
	 "001110000000000000001110",
	 "001110000000000000001110",
	 "001110000000000000011100",
	 "001110000000000000111000",
	 "001110000000000001110000",
	 "001110000000000111000000",
	 "001110000001110000000000",
	 "001110001111000000000000",
	 "001111111000000000000000"),
	 
	("001111111111111111111110",
	 "001111111111111111111110",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001111111111111111111110",
	 "001111111111111111111110",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001110000000000000000000",
	 "001111111111111111111110",
	 "001111111111111111111110"),
	 
	("000000000111100000000000",
	 "000000111000111000000000",
	 "000001110000001110000000",
	 "000111000000000011100000",
	 "001110000000000001110000",
	 "001110000000000001110000",
	 "001110000000000001110000",
	 "001111111111111111110000",
	 "001111111111111111110000",
	 "001110000000000001110000",
	 "001110000000000001110000",
	 "001110000000000001110000",
	 "001110000000000001110000",
	 "001110000000000001110000",
	 "001110000000000001110000"),
	 
	("001111110000000000000000",
	 "001111111110000000000000",
	 "001110000001110000000000",
	 "001110000000001110000000",
	 "001110000000000111100000",
	 "001110000000000000111000",
	 "001110000000000000001110",
	 "001110000000000000001110",
	 "001110000000000000011100",
	 "001110000000000000111000",
	 "001110000000000001110000",
	 "001110000000000111000000",
	 "001110000001110000000000",
	 "001110001111000000000000",
	 "001111111000000000000000"));
	  
	
	
end Num_Txt_Sprite;

package body Num_Txt_Sprite is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end Num_Txt_Sprite;
